// I2C TESTBENCH

module i2c_tb;
  reg clk,rst,newd,wr;
  reg [7:0] wdata;
  reg [6:0] addr;
  wire [7:0] rdata;
  wire done;
  
  i2c_design dut(clk,rst,newd,wr,wdata,addr,rdata,done);
  
  initial clk=0;
    always #5 clk=~clk;
  
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0,i2c_tb);
  end
  
  initial begin
    rst = 1;  //APPLY RESET
    newd = 0;
    wr = 0;
    wdata = 8'h00;
    addr = 7'h00;
    #20;
    rst = 0;  //RELEASE RESET
    #50;
      
    addr = 7'h10;
    wdata = $urandom_range(1,50); //8'h27;
    wr = 1'b1;
    newd = 1'b1;
    @(posedge done);  //WAIT FOR DONE SIGNAL
      
    newd = 1'b0;
    wr = 1'b0;
    #100;
      
    addr = 7'h10;
    wr = 1'b0;
    newd = 1'b1;
    @(posedge done);
    //if(rdata == 8'h27)
    if(wdata == rdata)
      $display("[PASS] : WDATA %0h -- %0h RDATA",wdata,rdata);
    else
      $display("[FAIL] : WDATA %0h -- %0h RDATA",wdata,rdata);
      
    #50;
    $finish();
    end
endmodule
